module iir_tb ();

localparam string in_file = "";
localparam string out_file = "";
localparam string cmp_file = "";

