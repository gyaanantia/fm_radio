`ifndef __GLOBALS__
`define __GLOBALS__

// UVM Globals
localparam string IQ_IN_NAME = "../read_iq.txt";
localparam string LEFT_OUT_NAME = "../left_out_uvm.txt";
localparam string RIGHT_OUT_NAME = "../right_out_uvm.txt";
localparam string RIGHT_CMP_NAME = "../right_volume.txt";
localparam string LEFT_CMP_NAME = "../left_volume.txt";
localparam int CLOCK_PERIOD = 10;

`endif
